entity ent is
END;

ARCHITECTURE arch OF ent IS
	 
BEGIN
END;

