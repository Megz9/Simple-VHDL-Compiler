entity ent is
END;

ARCHITECTURE arch OF ent IS
	SIGNAL s11 : t1;
	SIGNAL s11 : t1;
	SIGNAL s2 : t2;
BEGIN
	s11 <= s15;
	END;
